module alu32 (
    input [31:0] srca,
    input [31:0] srcb,
    input [3:0]  alucontrol,
    input [4:0]  shamt,
    output [31:0] aluout, 
    output zero);
);
    
endmodule